module ROM(a, out, clock);
input [8:0] a;
output reg [35:0] out;
reg [35:0] o;
input clock;
always @ (posedge clock)
begin
	out <= o;
end
always @(a) begin
case (a)
// --------- --- -- ------ --------- --- ----
// XXXXXXXXX JJJ SS FFEEII HOTCLSPMM WRF BBBB
// NEXT_ADDR MAA LR 01NNNN POPVPCVA REE 3210
// PMM LA ABVC CSP RR IAC
// CNZ 81 A TDT
// H
// --------- --- -- ------ --------- --- ----
9'h000 : o = 36'b000000010_000_00_000000_000000000_000_0000; // goto 0x2
9'h001 : o = 36'b001000000_000_00_110101_000000100_000_0001; // PC=PC+1;goto 0x40
9'h002 : o = 36'b000000000_100_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto (MBR)
9'h003 : o = 36'b000000100_000_00_010100_100000000_000_0111; // H=TOS;goto 0x4
9'h004 : o = 36'b000000010_000_00_111100_001000010_100_0000; // TOS=MDR=H+MDR;wr;goto 0x2
9'h005 : o = 36'b000000110_000_00_010100_100000000_000_0111; // H=TOS;goto 0x6
9'h006 : o = 36'b000000010_000_00_111111_001000010_100_0000; // TOS=MDR=MDR-H;wr;goto 0x2
9'h007 : o = 36'b000001000_000_00_010100_100000000_000_0111; // H=TOS;goto 0x8
9'h008 : o = 36'b000000010_000_00_001100_001000010_100_0000; // TOS=MDR=H AND MDR;wr;goto 0x2
9'h009 : o = 36'b000001010_000_00_010100_100000000_000_0111; // H=TOS;goto 0xA
9'h00a : o = 36'b000000010_000_00_011100_001000010_100_0000; // TOS=MDR=H OR MDR;wr;goto 0x2
9'h00b : o = 36'b000000010_000_00_010100_000000010_100_0111; // MDR=TOS;wr;goto 0x2
9'h00c : o = 36'b000001101_000_00_000000_000000000_000_0000; // goto 0xD
9'h00d : o = 36'b000000010_000_00_010100_001000000_000_0000; // TOS=MDR;goto 0x2
9'h00e : o = 36'b000001111_000_00_010100_000000001_000_0100; // MAR=SP;goto 0xF
9'h00f : o = 36'b000010001_000_00_010100_100000000_100_0000; // H=MDR;wr;goto 0x11
9'h010 : o = 36'b000010110_000_00_110101_000001001_000_0100; // SP=MAR=SP+1;goto 0x16
9'h011 : o = 36'b000010010_000_00_010100_000000010_000_0111; // MDR=TOS;goto 0x12
9'h012 : o = 36'b000010100_000_00_110110_000000001_100_0100; // MAR=SP-1;wr;goto 0x14
9'h013 : o = 36'b000100111_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x27
9'h014 : o = 36'b000000010_000_00_011000_001000000_000_0000; // TOS=H;goto 0x2
9'h015 : o = 36'b000011000_000_00_010100_100000000_000_0101; // H=LV;goto 0x18
9'h016 : o = 36'b000010111_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x17
9'h017 : o = 36'b000000010_000_00_010100_001000010_100_0010; // TOS=MDR=MBR;wr;goto 0x2
9'h018 : o = 36'b000011001_000_00_111100_000000001_010_0011; // MAR=H+MBRU;rd;goto 0x19
9'h019 : o = 36'b000011010_000_00_110101_000001001_000_0100; // SP=MAR=SP+1;goto 0x1A
9'h01a : o = 36'b000011011_000_00_110101_000000100_101_0001; // PC=PC+1;wr;fetch;goto 0x1B
9'h01b : o = 36'b000000010_000_00_010100_001000000_000_0000; // TOS=MDR;goto 0x2
9'h01c : o = 36'b000011101_000_00_111100_000000001_000_0011; // MAR=H+MBRU;goto 0x1D
9'h01d : o = 36'b000011110_000_00_010100_000000010_100_0111; // MDR=TOS;wr;goto 0x1E
9'h01e : o = 36'b000011111_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x1F
9'h01f : o = 36'b000100000_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x20
9'h020 : o = 36'b000000010_000_00_010100_001000000_000_0000; // TOS=MDR;goto 0x2
9'h021 : o = 36'b000100010_000_10_010100_100000000_000_0011; // H=MBRU<<8;goto 0x22
9'h022 : o = 36'b000100011_000_00_011100_100000000_000_0011; // H=H OR MBRU;goto 0x23
9'h023 : o = 36'b000011001_000_00_111100_000000001_010_0101; // MAR=H+LV;rd;goto 0x19
9'h024 : o = 36'b000100101_000_10_010100_100000000_000_0011; // H=MBRU<<8;goto 0x25
9'h025 : o = 36'b000100110_000_00_011100_100000000_000_0011; // H=H OR MBRU;goto 0x26
9'h026 : o = 36'b000011101_000_00_111100_000000001_000_0101; // MAR=H+LV;goto 0x1D
9'h027 : o = 36'b000101000_000_10_010100_100000000_000_0011; // H=MBRU<<8;goto 0x28
9'h028 : o = 36'b000101001_000_00_011100_100000000_000_0011; // H=H OR MBRU;goto 0x29
9'h029 : o = 36'b000011001_000_00_111100_000000001_010_0110; // MAR=H+CPP;rd;goto 0x19
9'h02a : o = 36'b000101011_000_00_111100_000000001_010_0011; // MAR=H+MBRU;rd;goto 0x2B
9'h02b : o = 36'b000101100_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x2C
9'h02c : o = 36'b000101101_000_00_010100_100000000_000_0000; // H=MDR;goto 0x2D
9'h02d : o = 36'b000101110_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x2E
9'h02e : o = 36'b000000010_000_00_111100_000000010_100_0010; // MDR=H+MBR;wr;goto 0x2
9'h02f : o = 36'b000110000_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x30
9'h030 : o = 36'b000110001_000_10_010100_100000000_000_0010; // H=MBR<<8;goto 0x31
9'h031 : o = 36'b000110010_000_00_011100_100000000_000_0011; // H=H OR MBRU;goto 0x32
9'h032 : o = 36'b000110011_000_00_111100_000000100_001_1000; // PC=H+OPC;fetch;goto 0x33
9'h033 : o = 36'b000000010_000_00_000000_000000000_000_0000; // goto 0x2
9'h034 : o = 36'b000110101_000_00_010100_010000000_000_0111; // OPC=TOS;goto 0x35
9'h035 : o = 36'b000110111_000_00_010100_001000000_000_0000; // TOS=MDR;goto 0x37
9'h036 : o = 36'b000011100_000_00_010100_100000000_000_0101; // H=LV;goto 0x1C
9'h037 : o = 36'b000000001_000_00_010100_000000000_000_1000; // N=OPC;if (N) goto 0x101; else goto 0x1
9'h038 : o = 36'b000111001_000_00_010100_010000000_000_0111; // OPC=TOS;goto 0x39
9'h039 : o = 36'b000111010_000_00_010100_001000000_000_0000; // TOS=MDR;goto 0x3A
9'h03a : o = 36'b000000001_011_00_010100_000000000_000_1000; // Z=OPC;if (Z) goto 0x101; else goto 0x1
9'h03b : o = 36'b000111100_000_00_110110_000001001_000_0100; // SP=MAR=SP-1;goto 0x3C
9'h03c : o = 36'b000111101_000_00_010100_100000000_010_0000; // H=MDR;rd;goto 0x3D
9'h03d : o = 36'b000111110_000_00_010100_010000000_000_0111; // OPC=TOS;goto 0x3E
9'h03e : o = 36'b000111111_000_00_010100_001000000_000_0000; // TOS=MDR;goto 0x3F
9'h03f : o = 36'b000000001_011_00_111111_000000000_000_1000; // Z=OPC-H;if (Z) goto 0x101; else goto 0x1
9'h040 : o = 36'b001000001_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x41
9'h041 : o = 36'b000000010_000_00_000000_000000000_000_0000; // goto 0x2
9'h042 : o = 36'b001000011_000_10_010100_100000000_000_0011; // H=MBRU<<8;goto 0x43
9'h043 : o = 36'b001000100_000_00_011100_100000000_000_0011; // H=H OR MBRU;goto 0x44
9'h044 : o = 36'b001000101_000_00_111100_000000001_010_0110; // MAR=H+CPP;rd;goto 0x45
9'h045 : o = 36'b001000110_000_00_110101_010000000_000_0001; // OPC=PC+1;goto 0x46
9'h046 : o = 36'b001000111_000_00_010100_000000100_001_0000; // PC=MDR;fetch;goto 0x47
9'h047 : o = 36'b001001000_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x48
9'h048 : o = 36'b001001001_000_10_010100_100000000_000_0011; // H=MBRU<<8;goto 0x49
9'h049 : o = 36'b001001010_000_00_011100_100000000_000_0011; // H=H OR MBRU;goto 0x4A
9'h04a : o = 36'b001001011_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x4B
9'h04b : o = 36'b001001100_000_00_111111_001000000_000_0100; // TOS=SP-H;goto 0x4C
9'h04c : o = 36'b001001101_000_00_110101_001000001_000_0111; // TOS=MAR=TOS+1;goto 0x4D
9'h04d : o = 36'b001001110_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x4E
9'h04e : o = 36'b001001111_000_10_010100_100000000_000_0011; // H=MBRU<<8;goto 0x4F
9'h04f : o = 36'b001010000_000_00_011100_100000000_000_0011; // H=H OR MBRU;goto 0x50
9'h050 : o = 36'b001010001_000_00_111101_000000010_100_0100; // MDR=H+SP+1;wr;goto 0x51
9'h051 : o = 36'b001010010_000_00_010100_000001001_000_0000; // SP=MAR=MDR;goto 0x52
9'h052 : o = 36'b001010011_000_00_010100_000000010_100_1000; // MDR=OPC;wr;goto 0x53
9'h053 : o = 36'b001010100_000_00_110101_000001001_000_0100; // SP=MAR=SP+1;goto 0x54
9'h054 : o = 36'b001010101_000_00_010100_000000010_100_0101; // MDR=LV;wr;goto 0x55
9'h055 : o = 36'b001010110_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x56
9'h056 : o = 36'b000000010_000_00_010100_000010000_000_0111; // LV=TOS;goto 0x2
9'h057 : o = 36'b000001100_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0xC
9'h058 : o = 36'b001011010_000_00_000000_000000000_000_0000; // goto 0x5A
9'h059 : o = 36'b000001011_000_00_110101_000001001_000_0100; // SP=MAR=SP+1;goto 0xB
9'h05a : o = 36'b001011011_000_00_010100_000010001_010_0000; // LV=MAR=MDR;rd;goto 0x5B
9'h05b : o = 36'b001011100_000_00_110101_000000001_000_0101; // MAR=LV+1;goto 0x5C
9'h05c : o = 36'b001011101_000_00_010100_000000100_011_0000; // PC=MDR;rd;fetch;goto 0x5D
9'h05d : o = 36'b001011110_000_00_010100_000000001_000_0100; // MAR=SP;goto 0x5E
9'h05e : o = 36'b001100001_000_00_010100_000010000_000_0000; // LV=MDR;goto 0x61
9'h05f : o = 36'b000001110_000_00_110110_000000001_010_0100; // MAR=SP-1;rd;goto 0xE
9'h060 : o = 36'b000000011_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x3
9'h061 : o = 36'b000000010_000_00_010100_000000010_100_0111; // MDR=TOS;wr;goto 0x2
9'h062 : o = 36'b001100011_000_00_010100_000000010_100_0111; // MDR=TOS;wr;goto 0x63
9'h063 : o = 36'b001100101_000_00_000000_000000000_000_0000; // goto 0x65
9'h064 : o = 36'b000000101_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x5
9'h065 : o = 36'b001100110_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x66
9'h066 : o = 36'b001100111_000_00_000000_000000000_000_0000; // goto 0x67
9'h067 : o = 36'b000000010_000_00_010100_001000000_000_0000; // TOS=MDR;goto 0x2
9'h068 : o = 36'b001101001_000_00_110101_000001001_000_0100; // SP=MAR=SP+1;goto 0x69
9'h069 : o = 36'b000000010_000_00_010100_001000000_100_0000; // TOS=MDR;wr;goto 0x2
9'h06a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h06b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h06c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h06d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h06e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h06f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h070 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h071 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h072 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h073 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h074 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h075 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h076 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h077 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h078 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h079 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h07a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h07b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h07c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h07d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h07e : o = 36'b000000111_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x7
9'h07f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h080 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h081 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h082 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h083 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h084 : o = 36'b000101010_000_00_010100_100000000_000_0101; // H=LV;goto 0x2A
9'h085 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h086 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h087 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h088 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h089 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h08a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h08b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h08c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h08d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h08e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h08f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h090 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h091 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h092 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h093 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h094 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h095 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h096 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h097 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h098 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h099 : o = 36'b000111000_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x38
9'h09a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h09b : o = 36'b000110100_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x34
9'h09c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h09d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h09e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h09f : o = 36'b000111011_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x3B
9'h0a0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a7 : o = 36'b000101111_000_00_110110_010000000_000_0001; // OPC=PC-1;goto 0x2F
9'h0a8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0a9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0aa : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ab : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ac : o = 36'b001011000_000_00_010100_000001001_010_0101; // SP=MAR=LV;rd;goto 0x58
9'h0ad : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ae : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0af : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b0 : o = 36'b000001001_000_00_110110_000001001_010_0100; // SP=MAR=SP-1;rd;goto 0x9
9'h0b1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b6 : o = 36'b001000010_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x42
9'h0b7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0b9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ba : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0bb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0bc : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0bd : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0be : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0bf : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c4 : o = 36'b100000000_100_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto (MBR OR 0x100)
9'h0c5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0c9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ca : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0cb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0cc : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0cd : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ce : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0cf : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0d9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0da : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0db : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0dc : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0dd : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0de : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0df : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0e9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ea : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0eb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ec : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ed : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ee : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ef : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0f9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0fa : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0fb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0fc : o = 36'b001101000_000_00_010010_000000001_010_0000; // MAR=-1;rd;goto 0x68
9'h0fd : o = 36'b001100010_000_00_010010_000000001_000_0000; // MAR=-1;goto 0x62
9'h0fe : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h0ff : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h100 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h101 : o = 36'b000101111_000_00_110110_010000000_001_0001; // OPC=PC-1;fetch;goto 0x2F
9'h102 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h103 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h104 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h105 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h106 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h107 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h108 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h109 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h10a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h10b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h10c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h10d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h10e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h10f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h110 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h111 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h112 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h113 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h114 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h115 : o = 36'b000100001_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x21
9'h116 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h117 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h118 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h119 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h11a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h11b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h11c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h11d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h11e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h11f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h120 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h121 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h122 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h123 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h124 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h125 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h126 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h127 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h128 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h129 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h12a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h12b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h12c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h12d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h12e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h12f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h130 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h131 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h132 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h133 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h134 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h135 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h136 : o = 36'b000100100_000_00_110101_000000100_001_0001; // PC=PC+1;fetch;goto 0x24
9'h137 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h138 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h139 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h13a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h13b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h13c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h13d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h13e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h13f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h140 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h141 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h142 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h143 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h144 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h145 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h146 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h147 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h148 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h149 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h14a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h14b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h14c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h14d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h14e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h14f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h150 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h151 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h152 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h153 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h154 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h155 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h156 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h157 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h158 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h159 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h15a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h15b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h15c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h15d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h15e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h15f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h160 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h161 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h162 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h163 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h164 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h165 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h166 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h167 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h168 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h169 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h16a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h16b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h16c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h16d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h16e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h16f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h170 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h171 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h172 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h173 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h174 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h175 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h176 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h177 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h178 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h179 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h17a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h17b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h17c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h17d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h17e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h17f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h180 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h181 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h182 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h183 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h184 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h185 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h186 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h187 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h188 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h189 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h18a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h18b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h18c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h18d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h18e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h18f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h190 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h191 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h192 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h193 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h194 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h195 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h196 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h197 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h198 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h199 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h19a : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h19b : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h19c : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h19d : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h19e : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h19f : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1a9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1aa : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ab : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ac : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ad : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ae : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1af : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1b9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ba : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1bb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1bc : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1bd : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1be : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1bf : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1c9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ca : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1cb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1cc : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1cd : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ce : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1cf : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1d9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1da : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1db : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1dc : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1dd : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1de : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1df : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1e9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ea : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1eb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ec : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ed : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ee : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ef : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f0 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f1 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f2 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f3 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f4 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f5 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f6 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f7 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f8 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1f9 : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1fa : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1fb : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1fc : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1fd : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1fe : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
9'h1ff : o = 36'b011111111_000_00_000000_000000000_000_0000; // goto 0xFF
endcase
end
endmodule